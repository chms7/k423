/*
 * @Design: k423_defines
 * @Author: Zhao Siwei 
 * @Email:  cheems@foxmail.com
 * @Date:   2023-11-11
 * @Description: Configuration of k423
 */

`define RST_PC 32'hFFFFFFFC
