/*
 * @Design: k423_if_bpu
 * @Author: Zhao Siwei 
 * @Email:  cheems@foxmail.com
 * @Date:   2023-12-10
 * @Description: Branch predict unit of if stage
 */
`include "k423_defines.svh"

module k423_if_bpu (
  // pc & instruction
  input logic [`CORE_ADDR_W -1:0] pc_i,
  input logic [`CORE_DATA_W -1:0] inst_i
);

endmodule
