/*
 * @Design: k423_defines
 * @Author: Zhao Siwei 
 * @Email:  cheems@foxmail.com
 * @Date:   2023-11-11
 * @Description: Configuration of k423
 */

// ---------------------------------------------------------------------------
// ISA
// ---------------------------------------------------------------------------
// `define ISA_M
`define ISA_Zicsr

// ---------------------------------------------------------------------------
// Reset PC
// ---------------------------------------------------------------------------
`define RST_PC      32'h0000_0000 - 32'd4

// ---------------------------------------------------------------------------
// Trap Base PC
// ---------------------------------------------------------------------------
`define TRAP_BASE   30'h00000000

// ---------------------------------------------------------------------------
// Branch Prediction
// ---------------------------------------------------------------------------
`define BPU_EN

// BHT
`define BHT_DEPTH   2
`define BHT_WIDTH   4

// PHT
`define PHT_DEPTH   32

// BTB
`define BTB_DEPTH   32

// RAS
`define RAS_DEPTH   8
